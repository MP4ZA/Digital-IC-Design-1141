module Mul_Mod (
    input  [22:0] A,
    input  [22:0] B,
    output [23:0] Z
);
/*
	Write Your Design Here ~
*/
    
endmodule
